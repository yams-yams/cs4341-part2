//-------------------------------------------------
//
// 4 to 16 decoder, Structural. 
// Group SAAMU Project Part 2
//
//-------------------------------------------------


//=================================================================
//
// DECODER
//
//=================================================================
module Dec(binary,onehot);

    input [3:0] binary;
    output [15:0]onehot;
    
    assign onehot[ 0]=~binary[3]&~binary[2]&~binary[1]&~binary[0];
    assign onehot[ 1]=~binary[3]&~binary[2]&~binary[1]& binary[0];
    assign onehot[ 2]=~binary[3]&~binary[2]& binary[1]&~binary[0];
    assign onehot[ 3]=~binary[3]&~binary[2]& binary[1]& binary[0];
    assign onehot[ 4]=~binary[3]& binary[2]&~binary[1]&~binary[0];
    assign onehot[ 5]=~binary[3]& binary[2]&~binary[1]& binary[0];
    assign onehot[ 6]=~binary[3]& binary[2]& binary[1]&~binary[0];
    assign onehot[ 7]=~binary[3]& binary[2]& binary[1]& binary[0];
    assign onehot[ 8]= binary[3]&~binary[2]&~binary[1]&~binary[0];
    assign onehot[ 9]= binary[3]&~binary[2]&~binary[1]& binary[0];
    assign onehot[10]= binary[3]&~binary[2]& binary[1]&~binary[0];
    assign onehot[11]= binary[3]&~binary[2]& binary[1]& binary[0];
    assign onehot[12]= binary[3]& binary[2]&~binary[1]&~binary[0];
    assign onehot[13]= binary[3]& binary[2]&~binary[1]& binary[0];
    assign onehot[14]= binary[3]& binary[2]& binary[1]&~binary[0];
    assign onehot[15]= binary[3]& binary[2]& binary[1]& binary[0];
	
endmodule
